magic
tech sky130A
magscale 1 2
timestamp 1729059214
<< error_s >>
rect 450 3483 456 3485
rect 719 3483 725 3485
rect 450 3479 725 3483
rect 444 3478 450 3479
rect 444 3473 448 3478
rect 725 3473 731 3479
rect 3507 3473 3706 3481
rect 3501 3467 3506 3473
rect 3708 3467 3712 3473
rect 444 3431 448 3437
rect 725 3431 731 3437
rect 3501 3431 3506 3435
rect 3708 3431 3712 3435
rect 450 3425 456 3431
rect 719 3425 725 3431
rect 3501 3429 3507 3431
rect 3706 3429 3712 3431
rect 3507 3423 3513 3429
rect 3700 3423 3706 3429
<< metal1 >>
rect 450 3922 3709 3971
rect 448 3431 450 3478
rect 863 3430 2045 3476
rect 2186 3431 3368 3477
rect 3506 3473 3708 3475
rect 3506 3431 3507 3473
rect 3706 3431 3708 3473
rect 450 2945 3709 2994
<< via1 >>
rect 450 3431 725 3479
rect 3507 3429 3706 3473
<< metal2 >>
rect 450 3922 3709 3971
rect 448 3431 450 3478
rect 3506 3473 3708 3475
rect 3506 3431 3507 3473
rect 3706 3431 3708 3473
rect 450 2945 3709 2994
use inverter2  x1
timestamp 1729055586
transform 1 0 848 0 1 4780
box -318 -1783 104 -857
use inverter2  x2
timestamp 1729055586
transform 1 0 2169 0 1 4780
box -318 -1783 104 -857
use inverter2  x3
timestamp 1729055586
transform 1 0 3490 0 1 4780
box -318 -1783 104 -857
<< end >>
