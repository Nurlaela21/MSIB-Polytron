magic
tech sky130A
magscale 1 2
timestamp 1729054860
<< viali >>
rect 918 -108 952 -32
rect 918 -638 952 -562
<< metal1 >>
rect 912 -32 958 -20
rect 912 -108 918 -32
rect 952 -108 1066 -32
rect 912 -120 958 -108
rect 1114 -120 1218 -86
rect 1076 -512 1110 -167
rect 1184 -550 1218 -120
rect 912 -562 958 -550
rect 912 -638 918 -562
rect 952 -638 1066 -562
rect 1114 -584 1218 -550
rect 912 -650 958 -638
use sky130_fd_pr__nfet_01v8_L9KS9E  XM1
timestamp 1729054860
transform 1 0 1093 0 1 -569
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_LJ7GBL  XM2
timestamp 1729054860
transform 1 0 1093 0 1 -106
box -211 -234 211 234
<< labels >>
flabel metal1 966 -88 1009 -52 0 FreeSans 160 0 0 0 VDD
port 1 nsew
flabel metal1 967 -615 1010 -579 0 FreeSans 160 0 0 0 GND
port 3 nsew
<< end >>
